library verilog;
use verilog.vl_types.all;
entity PROBLEM_3_vlg_vec_tst is
end PROBLEM_3_vlg_vec_tst;
