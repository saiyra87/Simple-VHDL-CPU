library verilog;
use verilog.vl_types.all;
entity PROBLEM_1_vlg_vec_tst is
end PROBLEM_1_vlg_vec_tst;
