library verilog;
use verilog.vl_types.all;
entity PROBLEM_2_vlg_vec_tst is
end PROBLEM_2_vlg_vec_tst;
